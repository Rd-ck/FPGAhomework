module FSM(
	input clk,
	input [3:0]b,
	output reg[3:0]a,
	output [7:0]seg);
reg[3:0] keyvalue;
reg[1:0] q=2'b0;

seg4_7 s0(
	.hex(keyvalue),
	.seg(seg)
	);

wire clk_4k;
clk_div #(1000) c0(
	.clk(clk),
	.clr(1),
	.clk_out(clk_4k)
	);
	
always @(posedge clk_4k)begin
	q<=q+1;
	case(q)
		0:a<=4'b1110;
		1:a<=4'b1101;
		2:a<=4'b1011;
		3:a<=4'b0111;
		default:a<=4'b0;
	endcase
	case ({a,b})
		8'b1110_0111: keyvalue<=4'h0;
		8'b1110_1011: keyvalue<=4'h1;
		8'b1110_1101: keyvalue<=4'h2;
		8'b1110_1110: keyvalue<=4'h3;
		
		8'b1101_0111: keyvalue<=4'h4;
		8'b1101_1011: keyvalue<=4'h5;
		8'b1101_1101: keyvalue<=4'h6;
		8'b1101_1110: keyvalue<=4'h7;
		
		8'b1011_0111: keyvalue<=4'h8;
		8'b1011_1011: keyvalue<=4'h9;
		8'b1011_1101: keyvalue<=4'ha;
		8'b1011_1110: keyvalue<=4'hb;
		
		8'b0111_0111: keyvalue<=4'hc;
		8'b0111_1011: keyvalue<=4'hd;
		8'b0111_1101: keyvalue<=4'he;
		8'b0111_1110: keyvalue<=4'hf;
	endcase
end

endmodule

