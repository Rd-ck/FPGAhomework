module fsm1_seq101(
	input clk,clr,x,
	output z);
	
reg [1:0]state;
parameter s0=2'b00,s1=2'b01,s2=2'b11,s3=2'b10;

always @(posedge clk or negedge clr)begin
	if(!clr)state <=s0;
	else begin
		case (state)
			s0:begin if(x) state<=s1;else state<=s0;end
			s1:begin if(x) state<=s1;else state<=s2;end
			s2:begin if(x) state<=s3;else state<=s0;end
			s3:begin if(x) state<=s1;else state<=s2;end
			default: state<=s0;
		endcase
	end
end

assign z=(state==s3)?1'b1:1'b0;

endmodule