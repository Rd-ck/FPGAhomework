module uart_rx
//========================< 参数 >==========================================
#(
parameter  CLK              = 50_000_000        , //系统时钟，50Mhz
parameter  BPS              = 9600              , //波特率
parameter  BPS_CNT          = CLK/BPS             //波特率计数
)
//========================< 端口 >==========================================
(
input   wire                clk                 , //时钟，50Mhz
input   wire                rst_n               , //复位，低电平有效
input   wire                din                 , //输入数据
output  reg   [7:0]         dout                , //输出数据
output  reg                 dout_vld              //输出数据的有效指示
);
//========================< 信号 >==========================================
reg                         rx0                 ;
reg                         rx1                 ;
reg                         rx2                 ;
wire                        rxv_en               ;
reg                         flag                ;
reg   [15:0]                cnt0                ;
wire                        add_cnt0            ;
wire                        end_cnt0            ;
reg   [ 3:0]                cnt1                ;
wire                        add_cnt1            ;
wire                        end_cnt1            ;
reg   [ 7:0]                data                ;

//==========================================================================
//==    消除亚稳态 + 下降沿检测
//==========================================================================
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        rx0 <= 1;
        rx1 <= 1;
        rx2 <= 1;
    end
    else begin
        rx0 <= din;
        rx1 <= rx0;
        rx2 <= rx1;
    end
end

assign rx_en = rx2 && ~rx1;

//==========================================================================
//==    接收状态指示
//==========================================================================
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        flag <= 0;
    else if(rx_en)
        flag <= 1;
    else if(end_cnt1)
        flag <= 0;
end

//==========================================================================
//==    波特率计数
//==========================================================================
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        cnt0 <= 0;
    else if(add_cnt0) begin
        if(end_cnt0)
            cnt0 <= 0;
        else
            cnt0 <= cnt0 + 1;
    end
end

assign add_cnt0 = flag;
assign end_cnt0 = cnt0== BPS_CNT-1 || end_cnt1;

//==========================================================================
//==    开始1位(不接收) + 数据8位 + 停止0.5位(不接收)，共10位
//==========================================================================
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        cnt1 <= 0;
    else if(add_cnt1) begin
        if(end_cnt1)
            cnt1 <= 0;
        else
            cnt1 <= cnt1 + 1;
    end
end

assign add_cnt1 = end_cnt0;
assign end_cnt1 = cnt1==10-1 && cnt0==BPS_CNT/2-1;

//==========================================================================
//==    缓存数据
//==========================================================================
always @ (posedge clk or negedge rst_n)begin
    if(!rst_n)
        data <= 8'd0;
    else if(cnt1>=1 && cnt1<=8 && cnt0==BPS_CNT/2-1) //中间采样
        data[cnt1-1] <= rx2;                         //或 dout <= {rx2,dout[7:1]};
end

//==========================================================================
//==    输出数据
//==========================================================================
always @ (posedge clk or negedge rst_n)begin
    if(!rst_n)
        dout <= 0;
    else if(end_cnt1)
        dout <= data;
end

always @ (posedge clk or negedge rst_n)begin
    if(!rst_n)
        dout_vld <= 0;
    else if(end_cnt1)
        dout_vld <= 1;
    else
        dout_vld <= 0;
end



endmodule